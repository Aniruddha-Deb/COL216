library ieee;
use ieee.std_logic_1164.all;

package Types is
    type signal_array is array(integer range <>) of std_logic_vector(integer range <>);

end Types;

package body MyTypes is
end MyTypes;
